version https://git-lfs.github.com/spec/v1
oid sha256:b495f453aad47999abcdbce5d2d47039b169e6c8ebcb7cd1e41ce2c0134c18f4
size 340241920

version https://git-lfs.github.com/spec/v1
oid sha256:a62d0a3672bbb255d43b8cd76b02f222c96ccbadaad260d8a46e650411d3d0a9
size 340241920

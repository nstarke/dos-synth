version https://git-lfs.github.com/spec/v1
oid sha256:43155bc05ee98a08c312b24d30f05030fa237a4e5b44bac1ce65b174c5eca2d9
size 340241920

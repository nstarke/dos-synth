version https://git-lfs.github.com/spec/v1
oid sha256:e45efa6f3301aaece43f67787670afe076c14426ffefd5baca25456b46d2de0a
size 340241920

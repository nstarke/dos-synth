version https://git-lfs.github.com/spec/v1
oid sha256:53eea50c9127bbb90d31cfa0cd60eab5d56961abab308f9c592c3cba8632a945
size 340241920
